module alu (A, B, FuncCode, C);

endmodule