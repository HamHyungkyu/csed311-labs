module register_file(read1, read2, write_reg, reg_write, write_data, read_out1, read_out2); 
    output read_out1;
    output read_out2;
    input read1;
    input read2;
    input reg_write;
    input write_reg;
    input write_data;
endmodule