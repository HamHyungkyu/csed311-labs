module register_file(read1, read2, write_reg, write_data, read_out1, read_out2); 
    output read_out1;
    output read_out2;
    input read1;
    input read2;
    input write_reg;
    input write_data;
endmodule